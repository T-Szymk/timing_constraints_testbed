// clocking block wrapper to contain instantiation of clocking wizard

module clock_wiz (
  input  logic clk,
  input  logic rst_n,   
  output logic clk_out  
  
);

endmodule : clock_wiz